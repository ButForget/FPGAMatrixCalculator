module transpose(input [3:0] a, output [3:0] o);


endmodule